module top_module ( input a, input b, output out );
    mod_a mod_a_0 (a, b, out);
endmodule